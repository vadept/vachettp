module vachettp_router

struct Controller_test {
}

pub fn (ct Controller_test) index() {}

fn test_route_from_path() {
	//GIVEN
	r := [
		Route{"path", Controller_test, "index"}
		]
	rtr := Router{r}

	//WHEN
	result = rtr.get_route_by_path ("path") or {}

	//THEN
	assert "path" == result.get_path()
	assert Controller_test == result.get_controller()
	assert "index" == result.get_method()
}

