module main

import vachettp

fn main() {
	vachettp.run_app()
}