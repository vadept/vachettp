module vachettp_router


